`include "src/const_param.v"

module mem_unit(
    input clk_in,
    input rst_in,
    input rdy_in,

    output wire mem_busy
);

endmodule
module instr_fetcher (
    
);
endmodule